
module frizzle;
endmodule
